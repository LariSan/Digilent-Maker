----------------------------------------------------------------------------------
-- Company: Digilent Romania
-- Engineer: Elod Gyorgy
-- 
-- Create Date:   11:44:47 01/12/2009
-- Modify Date:	06/03/2013
-- Design Name: 	
-- Module Name:  	Video - package
-- Project Name: 	Digilent VHDL Library
-- Target Devices: 
--
-- Tool versions: 
-- Description: This package defines video timing constants and the Digilent logo
-- bitmap.
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.04 - Added 1080P@60Hz
-- Revision 0.03 - Moved the Active Video area to the first part of the counter
-- Revision 0.02 - Added additional resolutions
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Video is


constant H_MAX : NATURAL := 4096;
constant V_MAX : NATURAL := 4096;
----------------------------------------------------------------------------------
-- Resolution selector enumeration
----------------------------------------------------------------------------------
type RESOLUTION is (R480_272P, R640_480P, R720_480P, R1280_720P, R1600_900P,
R800_600P, R800_480P, R1920_1080_60P, R1280_1024_60P, R1920_1080_30P);

----------------------------------------------------------------------------------
-- Timing Constants for 480x272 @60Hz
----------------------------------------------------------------------------------
--horizontal constants
constant H_480_272p_S : NATURAL := 45;		--sync
constant H_480_272p_FP : NATURAL := 0; 	--front porch
constant H_480_272p_AV : NATURAL := 480; 	--active video
constant H_480_272p_BP : NATURAL := 0;	--back porch
--vertical constants
constant V_480_272p_S : NATURAL := 16;		--sync
constant V_480_272p_FP : NATURAL := 0; 	--front porch
constant V_480_272p_AV : NATURAL := 272; 	--active video
constant V_480_272p_BP : NATURAL := 0;	--back porch

constant H_480_272p_AV_FP : NATURAL := H_480_272p_AV + H_480_272p_FP;
constant H_480_272p_AV_FP_S : NATURAL := H_480_272p_AV + H_480_272p_FP + H_480_272p_S;
constant H_480_272p_AV_FP_S_BP : NATURAL := H_480_272p_AV + H_480_272p_FP + H_480_272p_S + H_480_272p_BP;

constant V_480_272p_AV_FP : NATURAL := V_480_272p_AV + V_480_272p_FP;
constant V_480_272p_AV_FP_S : NATURAL := V_480_272p_AV + V_480_272p_FP + V_480_272p_S;
constant V_480_272p_AV_FP_S_BP : NATURAL := V_480_272p_AV + V_480_272p_FP + V_480_272p_S + V_480_272p_BP;

constant H_480_272p_POL : BOOLEAN := false; -- negative polarity
constant V_480_272p_POL : BOOLEAN := false; -- negative polarity

----------------------------------------------------------------------------------
-- Timing Constants for 640x480 @60Hz
----------------------------------------------------------------------------------
--horizontal constants
constant H_640_480p_S : NATURAL := 96;		--sync
constant H_640_480p_FP : NATURAL := 16; 	--front porch
constant H_640_480p_AV : NATURAL := 640; 	--active video
constant H_640_480p_BP : NATURAL := 48;	--back porch
--vertical constants
constant V_640_480p_S : NATURAL := 2;		--sync
constant V_640_480p_FP : NATURAL := 33; 	--front porch
constant V_640_480p_AV : NATURAL := 480; 	--active video
constant V_640_480p_BP : NATURAL := 10;	--back porch

constant H_640_480p_AV_FP : NATURAL := H_640_480p_AV + H_640_480p_FP;
constant H_640_480p_AV_FP_S : NATURAL := H_640_480p_AV + H_640_480p_FP + H_640_480p_S;
constant H_640_480p_AV_FP_S_BP : NATURAL := H_640_480p_AV + H_640_480p_FP + H_640_480p_S + H_640_480p_BP;

constant V_640_480p_AV_FP : NATURAL := V_640_480p_AV + V_640_480p_FP;
constant V_640_480p_AV_FP_S : NATURAL := V_640_480p_AV + V_640_480p_FP + V_640_480p_S;
constant V_640_480p_AV_FP_S_BP : NATURAL := V_640_480p_AV + V_640_480p_FP + V_640_480p_S + V_640_480p_BP;

constant H_640_480p_POL : BOOLEAN := false; -- negative polarity
constant V_640_480p_POL : BOOLEAN := false; -- negative polarity

----------------------------------------------------------------------------------
-- Timing Constants for 720x480 @60Hz
----------------------------------------------------------------------------------
--horizontal constants
constant H_720_480p_S : NATURAL := 62;		--sync
constant H_720_480p_FP : NATURAL := 16; 	--front porch
constant H_720_480p_AV : NATURAL := 720; 	--active video
constant H_720_480p_BP : NATURAL := 60;	--back porch
--vertical constants
constant V_720_480p_S : NATURAL := 6;		--sync
constant V_720_480p_FP : NATURAL := 9; 	--front porch
constant V_720_480p_AV : NATURAL := 480; 	--active video
constant V_720_480p_BP : NATURAL := 30;	--back porch

constant H_720_480p_AV_FP : NATURAL := H_720_480p_AV + H_720_480p_FP;
constant H_720_480p_AV_FP_S : NATURAL := H_720_480p_AV + H_720_480p_FP + H_720_480p_S;
constant H_720_480p_AV_FP_S_BP : NATURAL := H_720_480p_AV + H_720_480p_FP + H_720_480p_S + H_720_480p_BP;

constant V_720_480p_AV_FP : NATURAL := V_720_480p_AV + V_720_480p_FP;
constant V_720_480p_AV_FP_S : NATURAL := V_720_480p_AV + V_720_480p_FP + V_720_480p_S;
constant V_720_480p_AV_FP_S_BP : NATURAL := V_720_480p_AV + V_720_480p_FP + V_720_480p_S + V_720_480p_BP;

constant H_720_480p_POL : BOOLEAN := false; -- negative polarity
constant V_720_480p_POL : BOOLEAN := false; -- negative polarity

----------------------------------------------------------------------------------
-- Timing Constants for 1280x720 @60Hz 74.25MHz
----------------------------------------------------------------------------------
--horizontal constants
constant H_1280_720p_S : NATURAL := 40;		--sync
constant H_1280_720p_FP : NATURAL := 110; 	--front porch
constant H_1280_720p_AV : NATURAL := 1280; 	--active video
constant H_1280_720p_BP : NATURAL := 220;	--back porch
--vertical constants
constant V_1280_720p_S : NATURAL := 5;		--sync
constant V_1280_720p_FP : NATURAL := 5; 	--front porch
constant V_1280_720p_AV : NATURAL := 720; 	--active video
constant V_1280_720p_BP : NATURAL := 20;	--back porch

constant H_1280_720p_AV_FP : NATURAL := H_1280_720p_AV + H_1280_720p_FP;
constant H_1280_720p_AV_FP_S : NATURAL := H_1280_720p_AV + H_1280_720p_FP + H_1280_720p_S;
constant H_1280_720p_AV_FP_S_BP : NATURAL := H_1280_720p_AV + H_1280_720p_FP + H_1280_720p_S + H_1280_720p_BP;

constant V_1280_720p_AV_FP : NATURAL := V_1280_720p_AV + V_1280_720p_FP;
constant V_1280_720p_AV_FP_S : NATURAL := V_1280_720p_AV + V_1280_720p_FP + V_1280_720p_S;
constant V_1280_720p_AV_FP_S_BP : NATURAL := V_1280_720p_AV + V_1280_720p_FP + V_1280_720p_S + V_1280_720p_BP;

constant H_1280_720p_POL : BOOLEAN := true; -- positive polarity
constant V_1280_720p_POL : BOOLEAN := true; -- positive polarity

----------------------------------------------------------------------------------
-- Timing Constants for 1600x900 @60Hz 108MHz
----------------------------------------------------------------------------------
--horizontal constants
constant H_1600_900p_S : NATURAL := 20;		--sync
constant H_1600_900p_FP : NATURAL := 60; 	--front porch
constant H_1600_900p_AV : NATURAL := 1600; 	--active video
constant H_1600_900p_BP : NATURAL := 120;	--back porch
--vertical constants
constant V_1600_900p_S : NATURAL := 10;		--sync
constant V_1600_900p_FP : NATURAL := 20; 	--front porch
constant V_1600_900p_AV : NATURAL := 900; 	--active video
constant V_1600_900p_BP : NATURAL := 70;	--back porch

constant H_1600_900p_AV_FP : NATURAL := H_1600_900p_AV + H_1600_900p_FP;
constant H_1600_900p_AV_FP_S : NATURAL := H_1600_900p_AV + H_1600_900p_FP + H_1600_900p_S;
constant H_1600_900p_AV_FP_S_BP : NATURAL := H_1600_900p_AV + H_1600_900p_FP + H_1600_900p_S + H_1600_900p_BP;

constant V_1600_900p_AV_FP : NATURAL := V_1600_900p_AV + V_1600_900p_FP;
constant V_1600_900p_AV_FP_S : NATURAL := V_1600_900p_AV + V_1600_900p_FP + V_1600_900p_S;
constant V_1600_900p_AV_FP_S_BP : NATURAL := V_1600_900p_AV + V_1600_900p_FP + V_1600_900p_S + V_1600_900p_BP;

constant H_1600_900p_POL : BOOLEAN := true; -- positive polarity
constant V_1600_900p_POL : BOOLEAN := true; -- positive polarity

----------------------------------------------------------------------------------
-- Timing Constants for 800x600 @60Hz
----------------------------------------------------------------------------------
--horizontal constants
constant H_800_600p_S : NATURAL := 128;		--sync
constant H_800_600p_FP : NATURAL := 40; 	--front porch
constant H_800_600p_AV : NATURAL := 800; 	--active video
constant H_800_600p_BP : NATURAL := 88;	--back porch
--vertical constants
constant V_800_600p_S : NATURAL := 4;		--sync
constant V_800_600p_FP : NATURAL := 1; 	--front porch
constant V_800_600p_AV : NATURAL := 600; 	--active video
constant V_800_600p_BP : NATURAL := 23;	--back porch

constant H_800_600p_AV_FP : NATURAL := H_800_600p_AV + H_800_600p_FP;
constant H_800_600p_AV_FP_S : NATURAL := H_800_600p_AV + H_800_600p_FP + H_800_600p_S;
constant H_800_600p_AV_FP_S_BP : NATURAL := H_800_600p_AV + H_800_600p_FP + H_800_600p_S + H_800_600p_BP;

constant V_800_600p_AV_FP : NATURAL := V_800_600p_AV + V_800_600p_FP;
constant V_800_600p_AV_FP_S : NATURAL := V_800_600p_AV + V_800_600p_FP + V_800_600p_S;
constant V_800_600p_AV_FP_S_BP : NATURAL := V_800_600p_AV + V_800_600p_FP + V_800_600p_S + V_800_600p_BP;

constant H_800_600p_POL : BOOLEAN := true; -- positive polarity
constant V_800_600p_POL : BOOLEAN := true; -- positive polarity

----------------------------------------------------------------------------------
-- Timing Constants for 800x480 @60Hz
----------------------------------------------------------------------------------
--horizontal constants
constant H_800_480p_S : NATURAL := 1;		--sync
constant H_800_480p_FP : NATURAL := 1; 	--front porch
constant H_800_480p_AV : NATURAL := 800; 	--active video
constant H_800_480p_BP : NATURAL := 87;	--back porch
--vertical constants
constant V_800_480p_S : NATURAL := 3;		--sync
constant V_800_480p_FP : NATURAL := 1; 	--front porch
constant V_800_480p_AV : NATURAL := 480; 	--active video
constant V_800_480p_BP : NATURAL := 29;	--back porch

constant H_800_480p_AV_FP : NATURAL := H_800_480p_AV + H_800_480p_FP;
constant H_800_480p_AV_FP_S : NATURAL := H_800_480p_AV + H_800_480p_FP + H_800_480p_S;
constant H_800_480p_AV_FP_S_BP : NATURAL := H_800_480p_AV + H_800_480p_FP + H_800_480p_S + H_800_480p_BP;

constant V_800_480p_AV_FP : NATURAL := V_800_480p_AV + V_800_480p_FP;
constant V_800_480p_AV_FP_S : NATURAL := V_800_480p_AV + V_800_480p_FP + V_800_480p_S;
constant V_800_480p_AV_FP_S_BP : NATURAL := V_800_480p_AV + V_800_480p_FP + V_800_480p_S + V_800_480p_BP;

constant H_800_480p_POL : BOOLEAN := false; -- negative polarity
constant V_800_480p_POL : BOOLEAN := false; -- negative polarity

----------------------------------------------------------------------------------
-- Timing Constants for 1920x1080p @60Hz 148.5MHz
----------------------------------------------------------------------------------
--horizontal constants
constant H_1920_1080p_60_S : NATURAL := 44;		--sync
constant H_1920_1080p_60_FP : NATURAL := 88; 	--front porch
constant H_1920_1080p_60_AV : NATURAL := 1920; 	--active video
constant H_1920_1080p_60_BP : NATURAL := 148;	--back porch
--vertical constants
constant V_1920_1080p_60_S : NATURAL := 5;		--sync
constant V_1920_1080p_60_FP : NATURAL := 4; 	--front porch
constant V_1920_1080p_60_AV : NATURAL := 1080; 	--active video
constant V_1920_1080p_60_BP : NATURAL := 36;	--back porch

constant H_1920_1080p_60_AV_FP : NATURAL := H_1920_1080p_60_AV + H_1920_1080p_60_FP;
constant H_1920_1080p_60_AV_FP_S : NATURAL := H_1920_1080p_60_AV + H_1920_1080p_60_FP + H_1920_1080p_60_S;
constant H_1920_1080p_60_AV_FP_S_BP : NATURAL := H_1920_1080p_60_AV + H_1920_1080p_60_FP + H_1920_1080p_60_S + H_1920_1080p_60_BP;

constant V_1920_1080p_60_AV_FP : NATURAL := V_1920_1080p_60_AV + V_1920_1080p_60_FP;
constant V_1920_1080p_60_AV_FP_S : NATURAL := V_1920_1080p_60_AV + V_1920_1080p_60_FP + V_1920_1080p_60_S;
constant V_1920_1080p_60_AV_FP_S_BP : NATURAL := V_1920_1080p_60_AV + V_1920_1080p_60_FP + V_1920_1080p_60_S + V_1920_1080p_60_BP;

constant H_1920_1080p_60_POL : BOOLEAN := true; -- positive polarity
constant V_1920_1080p_60_POL : BOOLEAN := true; -- positive polarity

----------------------------------------------------------------------------------
-- Timing Constants for 1920x1080p @30Hz 74.25MHz
----------------------------------------------------------------------------------
--horizontal constants
constant H_1920_1080p_30_S : NATURAL := 44;		--sync
constant H_1920_1080p_30_FP : NATURAL := 88; 	--front porch
constant H_1920_1080p_30_AV : NATURAL := 1920; 	--active video
constant H_1920_1080p_30_BP : NATURAL := 148;	--back porch
--vertical constants
constant V_1920_1080p_30_S : NATURAL := 5;		--sync
constant V_1920_1080p_30_FP : NATURAL := 4; 	--front porch
constant V_1920_1080p_30_AV : NATURAL := 1080; 	--active video
constant V_1920_1080p_30_BP : NATURAL := 36;	--back porch

constant H_1920_1080p_30_AV_FP : NATURAL := H_1920_1080p_30_AV + H_1920_1080p_30_FP;
constant H_1920_1080p_30_AV_FP_S : NATURAL := H_1920_1080p_30_AV + H_1920_1080p_30_FP + H_1920_1080p_30_S;
constant H_1920_1080p_30_AV_FP_S_BP : NATURAL := H_1920_1080p_30_AV + H_1920_1080p_30_FP + H_1920_1080p_30_S + H_1920_1080p_30_BP;

constant V_1920_1080p_30_AV_FP : NATURAL := V_1920_1080p_30_AV + V_1920_1080p_30_FP;
constant V_1920_1080p_30_AV_FP_S : NATURAL := V_1920_1080p_30_AV + V_1920_1080p_30_FP + V_1920_1080p_30_S;
constant V_1920_1080p_30_AV_FP_S_BP : NATURAL := V_1920_1080p_30_AV + V_1920_1080p_30_FP + V_1920_1080p_30_S + V_1920_1080p_30_BP;

constant H_1920_1080p_30_POL : BOOLEAN := true; -- positive polarity
constant V_1920_1080p_30_POL : BOOLEAN := true; -- positive polarity

----------------------------------------------------------------------------------
-- Timing Constants for 1280x1024 @60Hz 108MHz
----------------------------------------------------------------------------------
--horizontal constants
constant H_1280_1024p_60_S : NATURAL := 112;		--sync
constant H_1280_1024p_60_FP : NATURAL := 48; 	--front porch
constant H_1280_1024p_60_AV : NATURAL := 1280; 	--active video
constant H_1280_1024p_60_BP : NATURAL := 248;	--back porch
--vertical constants
constant V_1280_1024p_60_S : NATURAL := 3;		--sync
constant V_1280_1024p_60_FP : NATURAL := 1; 	--front porch
constant V_1280_1024p_60_AV : NATURAL := 1024; 	--active video
constant V_1280_1024p_60_BP : NATURAL := 38;	--back porch

constant H_1280_1024p_60_AV_FP : NATURAL := H_1280_1024p_60_AV + H_1280_1024p_60_FP;
constant H_1280_1024p_60_AV_FP_S : NATURAL := H_1280_1024p_60_AV + H_1280_1024p_60_FP + H_1280_1024p_60_S;
constant H_1280_1024p_60_AV_FP_S_BP : NATURAL := H_1280_1024p_60_AV + H_1280_1024p_60_FP + H_1280_1024p_60_S + H_1280_1024p_60_BP;

constant V_1280_1024p_60_AV_FP : NATURAL := V_1280_1024p_60_AV + V_1280_1024p_60_FP;
constant V_1280_1024p_60_AV_FP_S : NATURAL := V_1280_1024p_60_AV + V_1280_1024p_60_FP + V_1280_1024p_60_S;
constant V_1280_1024p_60_AV_FP_S_BP : NATURAL := V_1280_1024p_60_AV + V_1280_1024p_60_FP + V_1280_1024p_60_S + V_1280_1024p_60_BP;

constant H_1280_1024p_60_POL : BOOLEAN := true; -- positive polarity
constant V_1280_1024p_60_POL : BOOLEAN := true; -- positive polarity

----------------------------------------------------------------------------------
-- Video ROM
----------------------------------------------------------------------------------
constant VROM_WIDTH : NATURAL := 250;
constant VROM_HEIGHT : NATURAL := 56;
constant VROM_COLOR_DEPTH : NATURAL := 16;
type vromt is array (0 to VROM_WIDTH*VROM_HEIGHT-1) of 
	std_logic_vector (VROM_COLOR_DEPTH-1 downto 0);
constant vrom : vromt := (
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"8430", x"528a", x"528a", x"528a", x"528a", x"528a", x"528a", x"7bcf", x"defb", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ce79", x"2104", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"1082", x"bdf7", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"2945", x"0000", x"0000", x"0000", x"2945", x"5acb", x"5acb", x"5acb", x"4a49", x"0882", x"0000", x"18c3", x"ef7d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"8c71", x"0000", x"0000", x"5acb", x"2945", x"738f", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"a534", x"18c3", x"0000", x"6b4d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"1082", x"0000", x"4a49", x"d6ba", x"b5b6", x"3186", x"b5b7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"7bcf", x"0000", x"0841", x"ce79", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5acb", x"0000", x"0841", x"bdf7", x"d6ba", x"d6ba", x"630c", x"738e", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"3186", x"0000", x"4208", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c638", x"0000", x"0000", x"6b8e", x"d6ba", x"d6ba", x"d6ba", x"c638", x"2945", x"ad76", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"9cf3", x"0000", x"0000", x"a534", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"3186", x"0000", x"2104", x"ce79", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8430", x"52cb", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"528a", x"0000", x"2104", x"ef7d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ce79", x"7bcf", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"4a49", x"0000", x"0000", x"94b2", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"3186", x"9cf4", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"ad75", x"1082", x"0000", x"4208", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"630c", x"7bcf", x"ce79", x"ffff", x"ffff", x"ffff",
x"ffff", x"f7be", x"630c", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"4208", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"a534", x"39c8", x"b5f7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"738e", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"6b4d", x"f7be", x"ffff",
x"ffff", x"6b4d", x"0000", x"0081", x"0245", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0943", x"0000", x"0841", x"b5b6", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4a49", x"8431", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"2945", x"0000", x"10c3", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0245", x"0081", x"0000", x"6b4d", x"ffff",
x"d6ba", x"0841", x"0081", x"0307", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"02c6", x"0000", x"0000", x"630c", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"bdf7", x"2945", x"b5b6", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"94b2", x"0000", x"0000", x"0286", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0081", x"0841", x"d6ba",
x"8c71", x"0000", x"0205", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0103", x"0000", x"18c3", x"ce79", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"6b4d", x"6b4d", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"4a49", x"0000", x"0882", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0205", x"0000", x"8c71",
x"630c", x"0000", x"0286", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0245", x"0000", x"0000", x"8c71", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce79", x"2945", x"ad75", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"ad75", x"1082", x"0000", x"0204", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"44ae", x"6d71", x"7db3", x"85f4", x"7db3", x"5d30", x"346c", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0388", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0387", x"0387", x"0387", x"0387", x"ffff", x"ffff", x"ffff", x"ffff", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0081", x"0000", x"3187", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8c71", x"8c71", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8c71", x"4a49", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"6b4d", x"0000", x"0041", x"0307", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"e77d", x"e77d", x"df7c", x"d73b", x"bef9", x"a676", x"7db3", x"3c6c", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"d73b", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"ae77", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"54ef", x"bef9", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e77d", x"9635", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"a676", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"df7c", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"5d30", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"346c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"a677", x"0387", x"0387", x"0387", x"0387", x"0387", x"85f4", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"e77d", x"2c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"e77d", x"13c9", x"0387", x"0387", x"0387", x"54ef", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"efbe", x"0b88", x"0387", x"0388", x"ffff", x"0388", x"0387", x"0387", x"0387", x"ffff", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"01c4", x"0000", x"0841", x"ad75", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"b5b7", x"0841", x"0841", x"bdf7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"39c7", x"94b3", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5b6", x"2104", x"0000", x"0943", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"df7c", x"6d71", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"3c6c", x"cf3a", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"8df4", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3b", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"5d2f", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"0b88", x"0b88", x"ffff", x"0387", x"ffff", x"ffff", x"ffff", x"0387", x"0387", x"ffff", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0040", x"0000", x"5acb", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4208", x"5acc", x"630c", x"4209", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"a535", x"3186", x"b5f7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"8c71", x"0000", x"0000", x"0ac6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3b", x"2c2b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"6531", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c6fa", x"1bca", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"5d2f", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"0b88", x"0b88", x"ffff", x"0387", x"ffff", x"0387", x"0387", x"ffff", x"0387", x"ffff", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0943", x"0000", x"1082", x"c638", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"94b2", x"3187", x"8cb2", x"94b2", x"39c7", x"9cf3", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"528a", x"7bcf", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"4208", x"0000", x"08c2", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbd", x"44ad", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"6d71", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"d73b", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"54ef", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"5d2f", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"0b88", x"0387", x"ffff", x"0387", x"ffff", x"ffff", x"ffff", x"0387", x"0387", x"ffff", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"0000", x"7c30", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce79", x"2945", x"7c30", x"94b2", x"94b2", x"8430", x"2945", x"ce7a", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"c638", x"2945", x"adb6", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"a534", x"0841", x"0000", x"0205", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbd", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"44ae", x"f7fe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbd", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"5d2f", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"0b88", x"0387", x"ffff", x"0387", x"ffff", x"0387", x"0387", x"ffff", x"0387", x"ffff", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"00c2", x"0000", x"2945", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"738e", x"4a4a", x"94b2", x"94b2", x"94b2", x"94b2", x"2946", x"738f", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"738e", x"630c", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"630c", x"0000", x"0041", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"85f4", x"6571", x"75b2", x"9635", x"c6fa", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"bef9", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"9635", x"3c6c", x"13c9", x"0b88", x"242b", x"7572", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"54ef", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"54ef", x"54ef", x"54ef", x"54ef", x"54ef", x"54ef", x"54ef", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c6f9", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"44ad", x"bef9", x"bef9", x"bef9", x"bef9", x"c6f9", x"f7ff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e77d", x"bef9", x"bef9", x"bef9", x"bef9", x"bef9", x"0b88", x"0387", x"0387", x"ffff", x"0387", x"0387", x"0387", x"0387", x"ffff", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0205", x"0000", x"0000", x"a534", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"bdf7", x"2104", x"8c71", x"94b2", x"94b2", x"94b2", x"94b2", x"3186", x"1082", x"bdf7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce79", x"2945", x"a534", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5b6", x"2104", x"0000", x"0984", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"2c2b", x"aeb8", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"44ae", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"75b2", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e77d", x"346c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"b6b8", x"ffff", x"ffff", x"c6fa", x"4cee", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"85f4", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ffff", x"ffff", x"ffff", x"ffff", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0041", x"0000", x"4a8a", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4a49", x"634d", x"94b2", x"94b2", x"94b2", x"94b2", x"8431", x"0841", x"0000", x"528a", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"94b2", x"4208", x"b5f7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"8430", x"0000", x"0000", x"0ac6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"a677", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"aeb8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7fe", x"3cad", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"9636", x"44ad", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"44ae", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0943", x"0000", x"1082", x"bdf7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"9cf3", x"3186", x"8cb2", x"94b2", x"94b2", x"94b2", x"94b2", x"39c7", x"0000", x"0000", x"0000", x"a534", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"39c8", x"8c72", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"39c7", x"0000", x"0102", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"efbd", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"346c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"a677", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e77d", x"13c9", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0ac6", x"0000", x"0000", x"738e", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce7a", x"2945", x"7bd0", x"94b2", x"94b2", x"94b2", x"94b2", x"738e", x"0000", x"0000", x"0841", x"0000", x"2945", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ad76", x"3186", x"b5b7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"9d34", x"0841", x"0000", x"0245", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"9e36", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"346c", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"6d71", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4cee", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"bef9", x"8df4", x"8df4", x"8df4", x"8df4", x"8df4", x"8df4", x"8df4", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e77d", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"aeb8", x"0388", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"08c2", x"0000", x"2104", x"ce7a", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"738e", x"4a49", x"94b2", x"94b2", x"94b2", x"94b2", x"8c72", x"2104", x"0000", x"0943", x"0286", x"0000", x"0000", x"8430", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"5acb", x"738e", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"5acb", x"0000", x"0081", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"6d71", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d2f", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"9635", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"13c9", x"0387", x"0387", x"0387", x"0387", x"2c2b", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"cf3a", x"9e36", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"44ad", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"6531", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"7572", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0205", x"0000", x"0000", x"9cf3", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"bdf7", x"2104", x"8c71", x"94b2", x"94b2", x"94b2", x"94b2", x"5acb", x"0000", x"0040", x"0307", x"0347", x"0943", x"0000", x"1082", x"c638", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"c638", x"2105", x"ad75", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"ad76", x"18c3", x"0000", x"01c4", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"a677", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbd", x"0388", x"0387", x"0387", x"0387", x"0387", x"346c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c6fa", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"44ad", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"a677", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"346c", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0041", x"0000", x"4208", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"528a", x"630c", x"94b2", x"94b2", x"94b2", x"94b2", x"8431", x"1082", x"0000", x"01c4", x"0387", x"0387", x"0307", x"0040", x"0000", x"5acb", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"7bcf", x"52cb", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"7bcf", x"0000", x"0000", x"0307", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"a677", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e77d", x"0388", x"0387", x"0387", x"0387", x"0387", x"346c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"bef9", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"44ad", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"13c9", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"d73b", x"13c9", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0984", x"0000", x"0841", x"b5f7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"a534", x"3186", x"8c72", x"94b2", x"94b2", x"94b2", x"8cb2", x"3a08", x"0000", x"0081", x"0347", x"0387", x"0387", x"0387", x"01c4", x"0000", x"0841", x"ad75", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ceba", x"3186", x"9cf4", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"3186", x"0000", x"0943", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"9635", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"0b88", x"0387", x"0387", x"0387", x"0387", x"346c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"aeb8", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"44ad", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"3c6c", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9e36", x"54ef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0ac6", x"0000", x"0000", x"6b4d", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"3186", x"7bcf", x"94b2", x"94b2", x"94b2", x"94b2", x"738f", x"0000", x"0000", x"0245", x"0387", x"0387", x"0387", x"0387", x"0347", x"0081", x"0000", x"3186", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"9cf3", x"39c7", x"b5f7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"94f3", x"0000", x"0000", x"0286", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"9635", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3cad", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"6d72", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242a", x"0387", x"0387", x"0387", x"0387", x"346c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c6fa", x"9e36", x"9e36", x"9e36", x"9e36", x"9e36", x"9e36", x"9e36", x"2c2b", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"7572", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"aeb8", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0102", x"0000", x"18c3", x"ce79", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"7bcf", x"4209", x"94b2", x"94b2", x"94b2", x"94b2", x"8c72", x"2104", x"0000", x"0102", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"0000", x"8c71", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4208", x"8430", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"528a", x"0000", x"0081", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"3c6c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6530", x"0387", x"0387", x"0387", x"0387", x"13c9", x"4cee", x"4cee", x"4cee", x"4cee", x"4cee", x"4cee", x"cf3a", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6531", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"b6b8", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0245", x"0000", x"0000", x"8c72", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"c638", x"2104", x"8c71", x"94b2", x"94b2", x"94b2", x"94b2", x"5acc", x"0000", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0103", x"0000", x"18c3", x"c679", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"b5b6", x"2945", x"b5b6", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"ad75", x"1082", x"0000", x"01c4", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"85f4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"bef9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c6fa", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"2c2b", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"1bc9", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0081", x"0000", x"39c7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"528a", x"5b0c", x"94b2", x"94b2", x"94b2", x"94b2", x"8431", x"1082", x"0000", x"0984", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0000", x"0000", x"630c", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"630c", x"6b4d", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"738e", x"0000", x"0041", x"0307", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"242b", x"0387", x"0387", x"0387", x"0387", x"13c9", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"85f4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d72", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"9635", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3b", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"44ad", x"f7fe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0984", x"0000", x"0841", x"b5b6", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"a535", x"2945", x"8c72", x"94b2", x"94b2", x"94b2", x"94b2", x"4208", x"0000", x"0041", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0984", x"0000", x"0841", x"b5b6", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce79", x"2145", x"a575", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5b7", x"2945", x"0000", x"0943", x"0347", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6d71", x"54ef", x"54ef", x"7572", x"a677", x"efbd", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3b", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"1bc9", x"e7bd", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"7572", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"9e36", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"6531", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"a676", x"85f4", x"85f4", x"85f4", x"85f4", x"85f4", x"85f4", x"85f4", x"346c", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"54ef", x"54ef", x"54ef", x"54ef", x"54ef", x"54ef", x"54ef", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"7db3", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0040", x"0000", x"5acc", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"3186", x"73cf", x"94b2", x"94b2", x"94b2", x"94b2", x"73cf", x"0000", x"0000", x"0245", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0041", x"0000", x"4208", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8430", x"4a4a", x"b5f7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"94b2", x"0000", x"0000", x"0ac6", x"0387", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"6531", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3b", x"7db3", x"54ef", x"44ae", x"6530", x"9635", x"e77d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3b", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"b6b8", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0103", x"0000", x"10c3", x"c638", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8430", x"4208", x"8cb2", x"94b2", x"94b2", x"94b2", x"8c72", x"2105", x"0000", x"08c2", x"0347", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0245", x"0000", x"0000", x"94b2", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"3186", x"94b3", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"4a49", x"0000", x"08c2", x"0347", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7fe", x"5d30", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"9e36", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"346c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"1bca", x"e77d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"0000", x"8430", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"c638", x"2104", x"8431", x"94b2", x"94b2", x"94b2", x"94b2", x"5acc", x"0000", x"0000", x"0ac6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"08c2", x"0000", x"2104", x"ce79", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"a534", x"3187", x"b5b7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"a575", x"1082", x"0000", x"0205", x"0387", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e7bd", x"4cee", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"9e36", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"4cee", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"4cee", x"f7fe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0081", x"0000", x"3186", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"5acb", x"5acb", x"94b2", x"94b2", x"94b2", x"94b2", x"8471", x"1082", x"0000", x"0984", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0ac6", x"0000", x"0000", x"6b8e", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4a4a", x"7bd0", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"6b4d", x"0000", x"0041", x"0307", x"0387", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"9e36", x"1bca", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"7572", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"d73b", x"3c6c", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"85f4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"02c6", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"01c4", x"0000", x"0000", x"a535", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ad75", x"2945", x"8c72", x"94b2", x"94b2", x"94b2", x"8cb2", x"4208", x"0000", x"0041", x"0307", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0984", x"0000", x"0841", x"bdf7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"bdf7", x"2104", x"b5b6", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5b6", x"2104", x"0000", x"0183", x"0347", x"0387", x"4cef", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"f7be", x"efbd", x"e77d", x"cf3a", x"a676", x"6530", x"1bc9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"df7c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"242a", x"9635", x"efbd", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"d73b", x"6d71", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"ae77", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"efbe", x"0b88", x"0387", x"0387", x"0387", x"0387", x"0387", x"6530", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5d30", x"0387", x"0387", x"0387", x"0b88", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b6b8", x"0387", x"0387", x"0387", x"0387", x"0387", x"8df4", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"cf3a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"c6f9", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"efbe", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9635", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"630c", x"0000", x"0286", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0040", x"0000", x"528a", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"39c7", x"738e", x"94b2", x"94b2", x"94b2", x"94b2", x"7bcf", x"0000", x"0000", x"0205", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0307", x"0041", x"0000", x"4a49", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"6b4d", x"630c", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"8c71", x"0000", x"0000", x"0ac6", x"0387", x"0b88", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"1bc9", x"1bc9", x"0b88", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"1bca", x"242a", x"242a", x"242a", x"242a", x"242a", x"1bc9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"44ae", x"7db3", x"9635", x"a677", x"ae77", x"a676", x"8df4", x"6531", x"2c2b", x"0388", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"1bc9", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"0b88", x"0387", x"0387", x"0387", x"0387", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"1bc9", x"0387", x"0387", x"0387", x"0387", x"0387", x"13c9", x"242a", x"242a", x"242a", x"242a", x"242a", x"1bca", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0b88", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"242a", x"242a", x"242a", x"242a", x"242a", x"242a", x"13c9", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0286", x"0000", x"738e",
x"8430", x"0000", x"0245", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"0943", x"0000", x"1082", x"c638", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8431", x"39c7", x"8cb2", x"94b2", x"94b2", x"94b2", x"8c72", x"2105", x"0000", x"0081", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0984", x"0000", x"0000", x"9cf3", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce79", x"2105", x"a534", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"4208", x"0000", x"08c2", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0245", x"0000", x"8430",
x"c638", x"0000", x"00c2", x"0347", x"0387", x"0387", x"0387", x"0387", x"0ac6", x"0000", x"0000", x"7bcf", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"c679", x"2104", x"8430", x"94b2", x"94b2", x"94b2", x"94b2", x"630c", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"18c3", x"a534", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4a49", x"4208", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"a534", x"0841", x"0000", x"0245", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0387", x"0347", x"00c2", x"0000", x"c638",
x"ffff", x"528a", x"0000", x"0103", x"0ac6", x"0347", x"0347", x"0b07", x"00c2", x"0000", x"2945", x"ce7a", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"630c", x"52cb", x"94b2", x"94b2", x"94b2", x"94b2", x"8c71", x"1082", x"0000", x"0841", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"1082", x"2945", x"3186", x"3186", x"3186", x"1082", x"3186", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"630c", x"0000", x"0081", x"0b07", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0ac6", x"0102", x"0000", x"528a", x"ffff",
x"ffff", x"ef7d", x"39c7", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"9cf3", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"b5b6", x"2105", x"8c72", x"94b2", x"94b2", x"94b2", x"94b2", x"4208", x"3186", x"9cf3", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5b6", x"18c3", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"4208", x"ef7d", x"ffff",
x"ffff", x"ffff", x"f7be", x"a534", x"528a", x"4208", x"3186", x"0000", x"0000", x"4a49", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4208", x"6b8e", x"94b2", x"94b2", x"94b2", x"94b2", x"7bcf", x"2104", x"adb6", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"8430", x"0000", x"0000", x"2945", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"4208", x"528a", x"a534", x"f7be", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5acb", x"0000", x"0841", x"bdf7", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"8c71", x"39c7", x"8cb2", x"94b2", x"94b2", x"94b2", x"8c72", x"2945", x"8430", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"b5f7", x"39c7", x"0000", x"4208", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c638", x"0000", x"0000", x"6b4d", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"ce79", x"2945", x"8430", x"94b2", x"94b2", x"94b2", x"94b2", x"630c", x"39c8", x"b5f7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"bdf7", x"9cf4", x"0841", x"0000", x"a534", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"d6ba", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"8430", x"b5b6", x"ffff", x"ffff", x"ffff", x"ffff", x"bdf7", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"bdf7", x"ffff", x"ce7a", x"7bd0", x"defb", x"ffff", x"ffff", x"ffff", x"b5b7", x"8430", x"ef7d", x"ffff", x"ffff", x"defb", x"7bcf", x"528a", x"4a49", x"738e", x"c679", x"ffff", x"ffff", x"ffff", x"ffff", x"defb", x"a575", x"ffff", x"ffff", x"ffff", x"f7be", x"8430", x"e73c", x"ffff", x"ffff", x"f7be", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"9cf3", x"e77d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"8c72", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"b5b6", x"ffff", x"f7be", x"8430", x"e73c", x"ffff", x"ffff", x"ffff", x"ffff", x"94f3", x"c638", x"ffff", x"ffff", x"ffff", x"94b2", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"ef7d", x"ffff", x"ffff", x"ffff", x"e73c", x"8430", x"528a", x"4a49", x"6b4d", x"bdf7", x"ffff", x"ffff", x"ffff", x"ffff", x"ef7d", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"7bd0", x"8c71", x"d6ba", x"ffff", x"ffff", x"ad75", x"8c71", x"f7be", x"ffff", x"ffff", x"ffff", x"94b2", x"9cf3", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5acb", x"0000", x"18c3", x"ce79", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"634d", x"528a", x"94b2", x"94b2", x"94b2", x"94b2", x"8c71", x"1082", x"630c", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"b5b6", x"ad75", x"1083", x"0000", x"39c7", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"1083", x"6b4e", x"6b4e", x"6b4e", x"630c", x"0882", x"ad75", x"ffff", x"ffff", x"ffff", x"8430", x"2104", x"6b4e", x"6b4e", x"6b4e", x"6b4e", x"6b4e", x"b5b6", x"ffff", x"f7be", x"630c", x"2945", x"e73c", x"ffff", x"bdf7", x"1082", x"9cf3", x"ffff", x"ffff", x"a575", x"1082", x"528b", x"94f3", x"9cf3", x"630c", x"1082", x"8430", x"ffff", x"ffff", x"ffff", x"c638", x"0841", x"a534", x"ffff", x"ffff", x"f7be", x"10c3", x"ce79", x"ffff", x"ffff", x"f7be", x"0841", x"5acb", x"6b4e", x"6b4d", x"39c7", x"18c3", x"c638", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"8c71", x"7bcf", x"7bcf", x"2104", x"4209", x"7bcf", x"7bcf", x"b5b6", x"ffff", x"e73c", x"0882", x"d6ba", x"ffff", x"ffff", x"ffff", x"ffff", x"39c7", x"94b2", x"ffff", x"ffff", x"ffff", x"31c7", x"4a49", x"6b4e", x"6b4e", x"6b4e", x"6b4e", x"6b4e", x"ef7d", x"ffff", x"ffff", x"bdf7", x"18c3", x"4a49", x"94b2", x"9d34", x"6b4d", x"1082", x"6b8e", x"ffff", x"ffff", x"ffff", x"d6fb", x"0841", x"630d", x"6b4e", x"6b4e", x"6b4e", x"4a8a", x"1082", x"defb", x"ffff", x"e73c", x"3186", x"630c", x"f7be", x"ffff", x"7bcf", x"2104", x"d6ba", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"3186", x"0000", x"4208", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"b5b7", x"2104", x"8c71", x"94b2", x"94b2", x"94b2", x"94b2", x"8430", x"2104", x"18c3", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"2104", x"18c3", x"0000", x"0000", x"1082", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"2145", x"ffff", x"ffff", x"ffff", x"ffff", x"39c7", x"8471", x"ffff", x"ffff", x"ffff", x"8430", x"4a49", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"5acb", x"3186", x"b5b6", x"10c3", x"94b2", x"ffff", x"ffff", x"e73c", x"1082", x"94b2", x"ffff", x"ffff", x"ffff", x"ffff", x"bdf7", x"0882", x"bdf7", x"ffff", x"ffff", x"c638", x"0841", x"1082", x"b5b6", x"ffff", x"f7be", x"10c3", x"ce79", x"ffff", x"ffff", x"f7be", x"0841", x"ceba", x"ffff", x"ffff", x"f7be", x"738e", x"2104", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4208", x"8c71", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"0882", x"d6ba", x"ffff", x"ffff", x"ffff", x"ffff", x"39c7", x"94b2", x"ffff", x"ffff", x"ffff", x"31c7", x"a534", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ef7d", x"2104", x"7c30", x"ffff", x"ffff", x"ffff", x"ffff", x"ce79", x"1083", x"a534", x"ffff", x"ffff", x"d6fb", x"0841", x"ef7d", x"ffff", x"ffff", x"ffff", x"f7be", x"18c4", x"ad75", x"ffff", x"ffff", x"defb", x"2145", x"6b4d", x"8431", x"18c3", x"ce79", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4a49", x"0000", x"2945", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"d6ba", x"4208", x"6b4d", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"8cb2", x"39c7", x"0000", x"2104", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"0882", x"39c7", x"39c7", x"39c7", x"3186", x"0882", x"d6ba", x"ffff", x"ffff", x"ffff", x"8430", x"18c4", x"528a", x"528a", x"528a", x"ad75", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"4a4a", x"0841", x"8c71", x"ffff", x"ffff", x"ffff", x"a534", x"2104", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4a49", x"738e", x"ffff", x"ffff", x"c638", x"2104", x"9cf3", x"1082", x"c638", x"f7be", x"10c3", x"ce79", x"ffff", x"ffff", x"f7be", x"0841", x"ceba", x"ffff", x"ffff", x"ffff", x"ef7d", x"0882", x"c638", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4208", x"8c71", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"0882", x"39c8", x"4a49", x"4a49", x"4a49", x"4a49", x"1083", x"94b2", x"ffff", x"ffff", x"ffff", x"31c7", x"39c7", x"528a", x"528a", x"528a", x"e73c", x"ffff", x"ffff", x"ffff", x"bdf7", x"1082", x"ef7d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"630d", x"5acb", x"ffff", x"ffff", x"d6fb", x"0841", x"738e", x"7bcf", x"7bcf", x"7bcf", x"5acb", x"1082", x"defb", x"ffff", x"ffff", x"ffff", x"d6ba", x"2104", x"18c3", x"c638", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"9cf3", x"0000", x"0000", x"94b2", x"d6ba", x"d6ba", x"d6ba", x"94b2", x"3186", x"8cb2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"8c72", x"18c3", x"0000", x"6b4d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"18c4", x"b5b6", x"b5b6", x"b5b6", x"ad75", x"528a", x"4a49", x"ffff", x"ffff", x"ffff", x"8430", x"2946", x"94f3", x"94f3", x"94f3", x"ce79", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"bdf7", x"10c3", x"f7be", x"ffff", x"ffff", x"ffff", x"9cf3", x"2945", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5acb", x"6b4d", x"ffff", x"ffff", x"c638", x"2104", x"f7be", x"8c71", x"18c3", x"c638", x"10c3", x"ce79", x"ffff", x"ffff", x"f7be", x"0841", x"ceba", x"ffff", x"ffff", x"ffff", x"ef7d", x"1082", x"bdf7", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4208", x"8c71", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"0882", x"8c71", x"a534", x"a534", x"a534", x"a534", x"2145", x"94b2", x"ffff", x"ffff", x"ffff", x"31c7", x"630c", x"94f3", x"94f3", x"94f3", x"ef7d", x"ffff", x"ffff", x"ffff", x"b5b6", x"18c3", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"738e", x"528b", x"ffff", x"ffff", x"d6fb", x"0841", x"634d", x"738e", x"738e", x"2945", x"2945", x"ce79", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"7bcf", x"5acb", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"f7be", x"3186", x"0000", x"2104", x"ce79", x"d6ba", x"ce79", x"2945", x"8430", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"528b", x"0000", x"1082", x"e73c", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"2145", x"ffff", x"ffff", x"ffff", x"ffff", x"c638", x"1082", x"ef7d", x"ffff", x"ffff", x"8430", x"4a49", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"be38", x"10c3", x"f7be", x"ffff", x"ffff", x"ffff", x"d6ba", x"0882", x"bdf7", x"ffff", x"ffff", x"ffff", x"ffff", x"defb", x"10c3", x"ad75", x"ffff", x"ffff", x"c638", x"2104", x"f7be", x"ffff", x"7bcf", x"18c4", x"0882", x"ce79", x"ffff", x"ffff", x"f7be", x"0841", x"ceba", x"ffff", x"ffff", x"ffff", x"a534", x"1082", x"ef7d", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4208", x"8c71", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"0882", x"d6ba", x"ffff", x"ffff", x"ffff", x"ffff", x"39c7", x"94b2", x"ffff", x"ffff", x"ffff", x"31c7", x"a534", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"1082", x"a534", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"2104", x"8cb2", x"ffff", x"ffff", x"d6fb", x"0841", x"ef7d", x"ffff", x"ffff", x"c638", x"1082", x"ce79", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"7c30", x"5acb", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"bdf7", x"0000", x"0000", x"738e", x"d6ba", x"6b4d", x"4a4a", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"8431", x"1082", x"0000", x"8c71", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"18c3", x"a534", x"a534", x"a534", x"a534", x"4a49", x"39c7", x"ffff", x"ffff", x"ffff", x"8430", x"3186", x"a534", x"a534", x"a534", x"a534", x"a534", x"b5f7", x"ffff", x"ffff", x"ffff", x"ffff", x"be38", x"10c3", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"7c30", x"10c3", x"8c71", x"ce79", x"ce79", x"9cf3", x"2104", x"528b", x"ffff", x"ffff", x"ffff", x"c638", x"2104", x"f7be", x"ffff", x"ffff", x"6b4d", x"0841", x"ce79", x"ffff", x"ffff", x"f7be", x"0841", x"8471", x"a534", x"9d34", x"6b4d", x"1082", x"94b2", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"4208", x"8c71", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"0882", x"d6ba", x"ffff", x"ffff", x"ffff", x"ffff", x"39c7", x"94b2", x"ffff", x"ffff", x"ffff", x"31c7", x"6b4d", x"a534", x"a534", x"a534", x"a534", x"a534", x"defb", x"ffff", x"ffff", x"94b2", x"1082", x"7bcf", x"c638", x"d6ba", x"a534", x"2945", x"4208", x"f7be", x"ffff", x"ffff", x"d6fb", x"0841", x"ef7d", x"ffff", x"ffff", x"ffff", x"73cf", x"39c7", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"7c30", x"5acb", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"5acb", x"0000", x"0841", x"4209", x"0841", x"8430", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"94b2", x"8471", x"3186", x"0000", x"2945", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"c638", x"4a49", x"4a49", x"4a49", x"4a49", x"4a49", x"6b8e", x"defb", x"ffff", x"ffff", x"ffff", x"a534", x"4a49", x"4a49", x"4a49", x"4a49", x"4a49", x"4a49", x"738e", x"ffff", x"ffff", x"ffff", x"ffff", x"ce79", x"528a", x"f7be", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ad75", x"4208", x"18c3", x"10c3", x"39c7", x"94b2", x"f7be", x"ffff", x"ffff", x"ffff", x"d6ba", x"5acb", x"f7be", x"ffff", x"ffff", x"f7be", x"738e", x"defb", x"ffff", x"ffff", x"f7be", x"4a49", x"4a49", x"4a49", x"4a49", x"6b4d", x"c638", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"738e", x"ad75", x"ffff", x"ffff", x"ffff", x"ffff", x"ef7d", x"4a49", x"defb", x"ffff", x"ffff", x"ffff", x"ffff", x"6b4d", x"ad76", x"ffff", x"ffff", x"ffff", x"6b4d", x"4a49", x"4a49", x"4a49", x"4a49", x"4a49", x"4a49", x"b5b6", x"ffff", x"ffff", x"ffff", x"bdf7", x"4a49", x"18c3", x"1083", x"3186", x"8c71", x"f7be", x"ffff", x"ffff", x"ffff", x"e73c", x"4a49", x"ef7d", x"ffff", x"ffff", x"ffff", x"ef7d", x"5acb", x"bdf7", x"ffff", x"ffff", x"ffff", x"ffff", x"a534", x"8430", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"defb", x"1082", x"0000", x"0000", x"0000", x"18c4", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"3186", x"1082", x"0000", x"0000", x"ad75", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"b5b6", x"18c3", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0841", x"94b2", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff",
x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"e73c", x"9cf3", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"7bcf", x"6b4d", x"8430", x"d6ba", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff", x"ffff");
attribute rom_extract : string;
attribute rom_style : string;
attribute rom_extract of vrom : constant is "yes";
attribute rom_style of vrom : constant is "block";
end Video;